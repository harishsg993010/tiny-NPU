// =============================================================================
// rsqrt_lut.sv - Inverse square root (1/sqrt(x)) approximation via 256-entry ROM
// Input:  x[15:0] unsigned (variance value, Q16.16 or raw unsigned)
// Output: rsqrt_out[15:0] unsigned (Q0.16 fixed-point)
// Index:  top 8 bits of x used as LUT index
// LUT:    rsqrt_lut[i] = round(65536 / sqrt(max(i,1) * 256))
//         i=0 special-cased to max value
// Pipeline: 1-cycle registered output
// =============================================================================
import npu_pkg::*;
import fixed_pkg::*;

module rsqrt_lut (
    input  logic        clk,
    input  logic [7:0]  addr,       // top 8 bits of variance
    output logic [15:0] data_out    // Q0.16 inverse square root
);

    // 256-entry ROM - inferred as block RAM
    (* rom_style = "block" *)
    logic [15:0] rom [0:255];

    // ----------------------------------------------------------------
    // ROM initialization
    // rsqrt_lut[i] = round(65536 / sqrt(i * 256))
    // = round(65536 / (16 * sqrt(i)))
    // = round(4096 / sqrt(i))
    // i=0 -> special: max value (65535)
    // i=1 -> 4096/1 = 4096
    // i=4 -> 4096/2 = 2048
    // i=16 -> 4096/4 = 1024
    // i=64 -> 4096/8 = 512
    // i=255 -> 4096/15.97 = 256
    // Placeholder values - regenerate with make_lut.py
    // ----------------------------------------------------------------
    initial begin
        rom[  0] = 16'hFFFF;  // special: 1/sqrt(0) = max
        rom[  1] = 16'd4096;  // 4096/sqrt(1)
        rom[  2] = 16'd2896;  // 4096/sqrt(2)
        rom[  3] = 16'd2365;  // 4096/sqrt(3)
        rom[  4] = 16'd2048;  // 4096/sqrt(4)
        rom[  5] = 16'd1832;
        rom[  6] = 16'd1672;
        rom[  7] = 16'd1548;
        rom[  8] = 16'd1448;
        rom[  9] = 16'd1365;
        rom[ 10] = 16'd1295;
        rom[ 11] = 16'd1235;
        rom[ 12] = 16'd1183;
        rom[ 13] = 16'd1136;
        rom[ 14] = 16'd1094;
        rom[ 15] = 16'd1058;
        rom[ 16] = 16'd1024;  // 4096/sqrt(16) = 1024
        rom[ 17] = 16'd993;
        rom[ 18] = 16'd966;
        rom[ 19] = 16'd940;
        rom[ 20] = 16'd916;
        rom[ 21] = 16'd894;
        rom[ 22] = 16'd873;
        rom[ 23] = 16'd854;
        rom[ 24] = 16'd836;
        rom[ 25] = 16'd819;   // 4096/sqrt(25) = 819
        rom[ 26] = 16'd803;
        rom[ 27] = 16'd788;
        rom[ 28] = 16'd774;
        rom[ 29] = 16'd761;
        rom[ 30] = 16'd748;
        rom[ 31] = 16'd736;
        rom[ 32] = 16'd724;
        rom[ 33] = 16'd713;
        rom[ 34] = 16'd702;
        rom[ 35] = 16'd692;
        rom[ 36] = 16'd683;   // 4096/sqrt(36) = 683
        rom[ 37] = 16'd673;
        rom[ 38] = 16'd664;
        rom[ 39] = 16'd656;
        rom[ 40] = 16'd648;
        rom[ 41] = 16'd640;
        rom[ 42] = 16'd632;
        rom[ 43] = 16'd625;
        rom[ 44] = 16'd617;
        rom[ 45] = 16'd611;
        rom[ 46] = 16'd604;
        rom[ 47] = 16'd597;
        rom[ 48] = 16'd591;
        rom[ 49] = 16'd585;   // 4096/sqrt(49) = 585
        rom[ 50] = 16'd579;
        rom[ 51] = 16'd573;
        rom[ 52] = 16'd568;
        rom[ 53] = 16'd563;
        rom[ 54] = 16'd557;
        rom[ 55] = 16'd552;
        rom[ 56] = 16'd547;
        rom[ 57] = 16'd543;
        rom[ 58] = 16'd538;
        rom[ 59] = 16'd533;
        rom[ 60] = 16'd529;
        rom[ 61] = 16'd524;
        rom[ 62] = 16'd520;
        rom[ 63] = 16'd516;
        rom[ 64] = 16'd512;   // 4096/sqrt(64) = 512
        rom[ 65] = 16'd508;
        rom[ 66] = 16'd504;
        rom[ 67] = 16'd500;
        rom[ 68] = 16'd497;
        rom[ 69] = 16'd493;
        rom[ 70] = 16'd489;
        rom[ 71] = 16'd486;
        rom[ 72] = 16'd483;
        rom[ 73] = 16'd479;
        rom[ 74] = 16'd476;
        rom[ 75] = 16'd473;
        rom[ 76] = 16'd470;
        rom[ 77] = 16'd467;
        rom[ 78] = 16'd464;
        rom[ 79] = 16'd461;
        rom[ 80] = 16'd458;
        rom[ 81] = 16'd455;   // 4096/sqrt(81) = 455
        rom[ 82] = 16'd452;
        rom[ 83] = 16'd450;
        rom[ 84] = 16'd447;
        rom[ 85] = 16'd444;
        rom[ 86] = 16'd442;
        rom[ 87] = 16'd439;
        rom[ 88] = 16'd437;
        rom[ 89] = 16'd434;
        rom[ 90] = 16'd432;
        rom[ 91] = 16'd429;
        rom[ 92] = 16'd427;
        rom[ 93] = 16'd425;
        rom[ 94] = 16'd422;
        rom[ 95] = 16'd420;
        rom[ 96] = 16'd418;
        rom[ 97] = 16'd416;
        rom[ 98] = 16'd414;
        rom[ 99] = 16'd411;
        rom[100] = 16'd410;   // 4096/sqrt(100) = 410
        rom[101] = 16'd408;
        rom[102] = 16'd406;
        rom[103] = 16'd404;
        rom[104] = 16'd402;
        rom[105] = 16'd400;
        rom[106] = 16'd398;
        rom[107] = 16'd396;
        rom[108] = 16'd394;
        rom[109] = 16'd392;
        rom[110] = 16'd390;
        rom[111] = 16'd389;
        rom[112] = 16'd387;
        rom[113] = 16'd385;
        rom[114] = 16'd384;
        rom[115] = 16'd382;
        rom[116] = 16'd380;
        rom[117] = 16'd379;
        rom[118] = 16'd377;
        rom[119] = 16'd375;
        rom[120] = 16'd374;
        rom[121] = 16'd372;   // 4096/sqrt(121) = 372
        rom[122] = 16'd371;
        rom[123] = 16'd369;
        rom[124] = 16'd368;
        rom[125] = 16'd366;
        rom[126] = 16'd365;
        rom[127] = 16'd363;
        rom[128] = 16'd362;
        rom[129] = 16'd360;
        rom[130] = 16'd359;
        rom[131] = 16'd358;
        rom[132] = 16'd356;
        rom[133] = 16'd355;
        rom[134] = 16'd354;
        rom[135] = 16'd352;
        rom[136] = 16'd351;
        rom[137] = 16'd350;
        rom[138] = 16'd348;
        rom[139] = 16'd347;
        rom[140] = 16'd346;
        rom[141] = 16'd345;
        rom[142] = 16'd343;
        rom[143] = 16'd342;
        rom[144] = 16'd341;   // 4096/sqrt(144) = 341
        rom[145] = 16'd340;
        rom[146] = 16'd339;
        rom[147] = 16'd338;
        rom[148] = 16'd337;
        rom[149] = 16'd335;
        rom[150] = 16'd334;
        rom[151] = 16'd333;
        rom[152] = 16'd332;
        rom[153] = 16'd331;
        rom[154] = 16'd330;
        rom[155] = 16'd329;
        rom[156] = 16'd328;
        rom[157] = 16'd327;
        rom[158] = 16'd326;
        rom[159] = 16'd325;
        rom[160] = 16'd324;
        rom[161] = 16'd323;
        rom[162] = 16'd322;
        rom[163] = 16'd321;
        rom[164] = 16'd320;
        rom[165] = 16'd319;
        rom[166] = 16'd318;
        rom[167] = 16'd317;
        rom[168] = 16'd316;
        rom[169] = 16'd315;   // 4096/sqrt(169) = 315
        rom[170] = 16'd314;
        rom[171] = 16'd313;
        rom[172] = 16'd312;
        rom[173] = 16'd311;
        rom[174] = 16'd311;
        rom[175] = 16'd310;
        rom[176] = 16'd309;
        rom[177] = 16'd308;
        rom[178] = 16'd307;
        rom[179] = 16'd306;
        rom[180] = 16'd305;
        rom[181] = 16'd305;
        rom[182] = 16'd304;
        rom[183] = 16'd303;
        rom[184] = 16'd302;
        rom[185] = 16'd301;
        rom[186] = 16'd300;
        rom[187] = 16'd300;
        rom[188] = 16'd299;
        rom[189] = 16'd298;
        rom[190] = 16'd297;
        rom[191] = 16'd296;
        rom[192] = 16'd296;
        rom[193] = 16'd295;
        rom[194] = 16'd294;
        rom[195] = 16'd293;
        rom[196] = 16'd293;   // 4096/sqrt(196) = 293
        rom[197] = 16'd292;
        rom[198] = 16'd291;
        rom[199] = 16'd291;
        rom[200] = 16'd290;
        rom[201] = 16'd289;
        rom[202] = 16'd288;
        rom[203] = 16'd288;
        rom[204] = 16'd287;
        rom[205] = 16'd286;
        rom[206] = 16'd286;
        rom[207] = 16'd285;
        rom[208] = 16'd284;
        rom[209] = 16'd284;
        rom[210] = 16'd283;
        rom[211] = 16'd282;
        rom[212] = 16'd282;
        rom[213] = 16'd281;
        rom[214] = 16'd280;
        rom[215] = 16'd280;
        rom[216] = 16'd279;
        rom[217] = 16'd278;
        rom[218] = 16'd278;
        rom[219] = 16'd277;
        rom[220] = 16'd276;
        rom[221] = 16'd276;
        rom[222] = 16'd275;
        rom[223] = 16'd275;
        rom[224] = 16'd274;
        rom[225] = 16'd273;   // 4096/sqrt(225) = 273
        rom[226] = 16'd273;
        rom[227] = 16'd272;
        rom[228] = 16'd271;
        rom[229] = 16'd271;
        rom[230] = 16'd270;
        rom[231] = 16'd270;
        rom[232] = 16'd269;
        rom[233] = 16'd268;
        rom[234] = 16'd268;
        rom[235] = 16'd267;
        rom[236] = 16'd267;
        rom[237] = 16'd266;
        rom[238] = 16'd266;
        rom[239] = 16'd265;
        rom[240] = 16'd264;
        rom[241] = 16'd264;
        rom[242] = 16'd263;
        rom[243] = 16'd263;
        rom[244] = 16'd262;
        rom[245] = 16'd262;
        rom[246] = 16'd261;
        rom[247] = 16'd261;
        rom[248] = 16'd260;
        rom[249] = 16'd260;
        rom[250] = 16'd259;
        rom[251] = 16'd259;
        rom[252] = 16'd258;
        rom[253] = 16'd258;
        rom[254] = 16'd257;
        rom[255] = 16'd256;   // 4096/sqrt(255) ~ 257
    end

    // ----------------------------------------------------------------
    // Registered read (1-cycle latency)
    // ----------------------------------------------------------------
    always_ff @(posedge clk) begin
        data_out <= rom[addr];
    end

endmodule
