// =============================================================================
// graph_exp_lut.sv - EXP activation function via 256-entry ROM lookup table
// Input:  x[7:0] signed int8
// Output: data_out[7:0] signed int8
// Formula: LUT[i] = clamp(round(exp(signed_i / 32) * 32), -128, 127)
// Scale: int8 maps to float via /32, so int8 range [-128,127] -> [-4.0, 3.97]
// Pipeline: 1-cycle registered output
// =============================================================================
`default_nettype none

module graph_exp_lut (
    input  wire        clk,
    input  wire  [7:0] addr,       // treated as signed int8 index
    output logic [7:0] data_out    // signed int8 EXP result
);

    // 256-entry ROM - inferred as block RAM
    (* rom_style = "block" *)
    logic [7:0] rom [0:255];

    // ----------------------------------------------------------------
    // ROM initialization
    // LUT[i] = clamp(round(exp(signed_i / 32.0) * 32.0), -128, 127)
    //
    // Key values (signed int8 index -> EXP output):
    //   0   -> 32  (exp(0)*32 = 32)
    //   32  -> 87  (exp(1)*32 = 86.99)
    //   64  -> 127 (exp(2)*32 = 236.4 -> clamped)
    //  -32  -> 12  (exp(-1)*32 = 11.77)
    //  -128 -> 1   (exp(-4)*32 = 0.586)
    // ----------------------------------------------------------------
    initial begin
        // Positive indices 0..127 (signed 0 to +127)
        // x_float = i/32.0, range [0, 3.97]
        rom[  0] = 8'h20;    // exp(0.000)*32 = 32
        rom[  1] = 8'h21;    // 33
        rom[  2] = 8'h22;    // 34
        rom[  3] = 8'h23;    // 35
        rom[  4] = 8'h24;    // 36
        rom[  5] = 8'h25;    // 37
        rom[  6] = 8'h27;    // 39
        rom[  7] = 8'h28;    // 40
        rom[  8] = 8'h29;    // 41
        rom[  9] = 8'h2A;    // 42
        rom[ 10] = 8'h2C;    // 44
        rom[ 11] = 8'h2D;    // 45
        rom[ 12] = 8'h2F;    // 47
        rom[ 13] = 8'h30;    // 48
        rom[ 14] = 8'h32;    // 50
        rom[ 15] = 8'h33;    // 51
        rom[ 16] = 8'h35;    // 53  exp(0.5)*32
        rom[ 17] = 8'h36;    // 54
        rom[ 18] = 8'h38;    // 56
        rom[ 19] = 8'h3A;    // 58
        rom[ 20] = 8'h3C;    // 60
        rom[ 21] = 8'h3E;    // 62
        rom[ 22] = 8'h40;    // 64
        rom[ 23] = 8'h42;    // 66
        rom[ 24] = 8'h44;    // 68
        rom[ 25] = 8'h46;    // 70
        rom[ 26] = 8'h48;    // 72
        rom[ 27] = 8'h4A;    // 74
        rom[ 28] = 8'h4D;    // 77
        rom[ 29] = 8'h4F;    // 79
        rom[ 30] = 8'h52;    // 82
        rom[ 31] = 8'h54;    // 84
        rom[ 32] = 8'h57;    // 87  exp(1.0)*32
        rom[ 33] = 8'h5A;    // 90
        rom[ 34] = 8'h5D;    // 93
        rom[ 35] = 8'h60;    // 96
        rom[ 36] = 8'h63;    // 99
        rom[ 37] = 8'h66;    // 102
        rom[ 38] = 8'h69;    // 105
        rom[ 39] = 8'h6C;    // 108
        rom[ 40] = 8'h70;    // 112
        rom[ 41] = 8'h73;    // 115
        rom[ 42] = 8'h77;    // 119
        rom[ 43] = 8'h7B;    // 123
        rom[ 44] = 8'h7F;    // 127 (clamped)
        rom[ 45] = 8'h7F;    // 127
        rom[ 46] = 8'h7F;    // 127
        rom[ 47] = 8'h7F;    // 127
        rom[ 48] = 8'h7F;    // 127  exp(1.5)*32 = 143 -> clamped
        rom[ 49] = 8'h7F;
        rom[ 50] = 8'h7F;
        rom[ 51] = 8'h7F;
        rom[ 52] = 8'h7F;
        rom[ 53] = 8'h7F;
        rom[ 54] = 8'h7F;
        rom[ 55] = 8'h7F;
        rom[ 56] = 8'h7F;
        rom[ 57] = 8'h7F;
        rom[ 58] = 8'h7F;
        rom[ 59] = 8'h7F;
        rom[ 60] = 8'h7F;
        rom[ 61] = 8'h7F;
        rom[ 62] = 8'h7F;
        rom[ 63] = 8'h7F;
        rom[ 64] = 8'h7F;    // exp(2.0)*32 = 236 -> clamped
        rom[ 65] = 8'h7F;
        rom[ 66] = 8'h7F;
        rom[ 67] = 8'h7F;
        rom[ 68] = 8'h7F;
        rom[ 69] = 8'h7F;
        rom[ 70] = 8'h7F;
        rom[ 71] = 8'h7F;
        rom[ 72] = 8'h7F;
        rom[ 73] = 8'h7F;
        rom[ 74] = 8'h7F;
        rom[ 75] = 8'h7F;
        rom[ 76] = 8'h7F;
        rom[ 77] = 8'h7F;
        rom[ 78] = 8'h7F;
        rom[ 79] = 8'h7F;
        rom[ 80] = 8'h7F;
        rom[ 81] = 8'h7F;
        rom[ 82] = 8'h7F;
        rom[ 83] = 8'h7F;
        rom[ 84] = 8'h7F;
        rom[ 85] = 8'h7F;
        rom[ 86] = 8'h7F;
        rom[ 87] = 8'h7F;
        rom[ 88] = 8'h7F;
        rom[ 89] = 8'h7F;
        rom[ 90] = 8'h7F;
        rom[ 91] = 8'h7F;
        rom[ 92] = 8'h7F;
        rom[ 93] = 8'h7F;
        rom[ 94] = 8'h7F;
        rom[ 95] = 8'h7F;
        rom[ 96] = 8'h7F;    // exp(3.0)*32 = 643 -> clamped
        rom[ 97] = 8'h7F;
        rom[ 98] = 8'h7F;
        rom[ 99] = 8'h7F;
        rom[100] = 8'h7F;
        rom[101] = 8'h7F;
        rom[102] = 8'h7F;
        rom[103] = 8'h7F;
        rom[104] = 8'h7F;
        rom[105] = 8'h7F;
        rom[106] = 8'h7F;
        rom[107] = 8'h7F;
        rom[108] = 8'h7F;
        rom[109] = 8'h7F;
        rom[110] = 8'h7F;
        rom[111] = 8'h7F;
        rom[112] = 8'h7F;
        rom[113] = 8'h7F;
        rom[114] = 8'h7F;
        rom[115] = 8'h7F;
        rom[116] = 8'h7F;
        rom[117] = 8'h7F;
        rom[118] = 8'h7F;
        rom[119] = 8'h7F;
        rom[120] = 8'h7F;
        rom[121] = 8'h7F;
        rom[122] = 8'h7F;
        rom[123] = 8'h7F;
        rom[124] = 8'h7F;
        rom[125] = 8'h7F;
        rom[126] = 8'h7F;
        rom[127] = 8'h7F;

        // Negative indices 128..255 (signed -128 to -1)
        // x_float = (i-256)/32.0, range [-4.0, -0.03125]
        // exp() of negative values -> small positive results
        rom[128] = 8'h01;    // exp(-4.000)*32 = 0.59 -> 1
        rom[129] = 8'h01;    // exp(-3.969)*32 = 0.60
        rom[130] = 8'h01;    // exp(-3.938)*32 = 0.62
        rom[131] = 8'h01;    // exp(-3.906)*32 = 0.64
        rom[132] = 8'h01;    // exp(-3.875)*32 = 0.66
        rom[133] = 8'h01;    // exp(-3.844)*32 = 0.69
        rom[134] = 8'h01;    // exp(-3.813)*32 = 0.71
        rom[135] = 8'h01;    // exp(-3.781)*32 = 0.73
        rom[136] = 8'h01;    // exp(-3.750)*32 = 0.75
        rom[137] = 8'h01;    // exp(-3.719)*32 = 0.78
        rom[138] = 8'h01;    // exp(-3.688)*32 = 0.80
        rom[139] = 8'h01;    // exp(-3.656)*32 = 0.83
        rom[140] = 8'h01;    // exp(-3.625)*32 = 0.85
        rom[141] = 8'h01;    // exp(-3.594)*32 = 0.88
        rom[142] = 8'h01;    // exp(-3.563)*32 = 0.91
        rom[143] = 8'h01;    // exp(-3.531)*32 = 0.94
        rom[144] = 8'h01;    // exp(-3.500)*32 = 0.97 -> 1
        rom[145] = 8'h01;    // exp(-3.469)*32 = 1.00
        rom[146] = 8'h01;    // exp(-3.438)*32 = 1.03
        rom[147] = 8'h01;    // exp(-3.406)*32 = 1.06
        rom[148] = 8'h01;    // exp(-3.375)*32 = 1.10
        rom[149] = 8'h01;    // exp(-3.344)*32 = 1.13
        rom[150] = 8'h01;    // exp(-3.313)*32 = 1.17
        rom[151] = 8'h01;    // exp(-3.281)*32 = 1.20
        rom[152] = 8'h01;    // exp(-3.250)*32 = 1.24
        rom[153] = 8'h01;    // exp(-3.219)*32 = 1.28
        rom[154] = 8'h01;    // exp(-3.188)*32 = 1.32
        rom[155] = 8'h01;    // exp(-3.156)*32 = 1.36
        rom[156] = 8'h01;    // exp(-3.125)*32 = 1.41
        rom[157] = 8'h01;    // exp(-3.094)*32 = 1.45
        rom[158] = 8'h01;    // exp(-3.063)*32 = 1.50
        rom[159] = 8'h02;    // exp(-3.031)*32 = 1.55 -> 2
        rom[160] = 8'h02;    // exp(-3.000)*32 = 1.59 -> 2
        rom[161] = 8'h02;    // exp(-2.969)*32 = 1.64
        rom[162] = 8'h02;    // exp(-2.938)*32 = 1.70
        rom[163] = 8'h02;    // exp(-2.906)*32 = 1.75
        rom[164] = 8'h02;    // exp(-2.875)*32 = 1.81
        rom[165] = 8'h02;    // exp(-2.844)*32 = 1.86
        rom[166] = 8'h02;    // exp(-2.813)*32 = 1.92
        rom[167] = 8'h02;    // exp(-2.781)*32 = 1.98
        rom[168] = 8'h02;    // exp(-2.750)*32 = 2.05
        rom[169] = 8'h02;    // exp(-2.719)*32 = 2.11
        rom[170] = 8'h02;    // exp(-2.688)*32 = 2.18
        rom[171] = 8'h02;    // exp(-2.656)*32 = 2.25
        rom[172] = 8'h02;    // exp(-2.625)*32 = 2.32
        rom[173] = 8'h02;    // exp(-2.594)*32 = 2.39
        rom[174] = 8'h02;    // exp(-2.563)*32 = 2.47
        rom[175] = 8'h03;    // exp(-2.531)*32 = 2.55 -> 3
        rom[176] = 8'h03;    // exp(-2.500)*32 = 2.63 -> 3
        rom[177] = 8'h03;    // exp(-2.469)*32 = 2.71
        rom[178] = 8'h03;    // exp(-2.438)*32 = 2.80
        rom[179] = 8'h03;    // exp(-2.406)*32 = 2.89
        rom[180] = 8'h03;    // exp(-2.375)*32 = 2.98
        rom[181] = 8'h03;    // exp(-2.344)*32 = 3.07
        rom[182] = 8'h03;    // exp(-2.313)*32 = 3.17
        rom[183] = 8'h03;    // exp(-2.281)*32 = 3.27
        rom[184] = 8'h03;    // exp(-2.250)*32 = 3.37
        rom[185] = 8'h03;    // exp(-2.219)*32 = 3.48
        rom[186] = 8'h04;    // exp(-2.188)*32 = 3.59 -> 4
        rom[187] = 8'h04;    // exp(-2.156)*32 = 3.71
        rom[188] = 8'h04;    // exp(-2.125)*32 = 3.83
        rom[189] = 8'h04;    // exp(-2.094)*32 = 3.95
        rom[190] = 8'h04;    // exp(-2.063)*32 = 4.07
        rom[191] = 8'h04;    // exp(-2.031)*32 = 4.20
        rom[192] = 8'h04;    // exp(-2.000)*32 = 4.33 -> 4
        rom[193] = 8'h04;    // exp(-1.969)*32 = 4.47
        rom[194] = 8'h05;    // exp(-1.938)*32 = 4.61 -> 5
        rom[195] = 8'h05;    // exp(-1.906)*32 = 4.76
        rom[196] = 8'h05;    // exp(-1.875)*32 = 4.91
        rom[197] = 8'h05;    // exp(-1.844)*32 = 5.07
        rom[198] = 8'h05;    // exp(-1.813)*32 = 5.23
        rom[199] = 8'h05;    // exp(-1.781)*32 = 5.39
        rom[200] = 8'h06;    // exp(-1.750)*32 = 5.57 -> 6
        rom[201] = 8'h06;    // exp(-1.719)*32 = 5.75
        rom[202] = 8'h06;    // exp(-1.688)*32 = 5.93
        rom[203] = 8'h06;    // exp(-1.656)*32 = 6.12
        rom[204] = 8'h06;    // exp(-1.625)*32 = 6.32
        rom[205] = 8'h07;    // exp(-1.594)*32 = 6.52 -> 7
        rom[206] = 8'h07;    // exp(-1.563)*32 = 6.73
        rom[207] = 8'h07;    // exp(-1.531)*32 = 6.95
        rom[208] = 8'h07;    // exp(-1.500)*32 = 7.14 -> 7
        rom[209] = 8'h07;    // exp(-1.469)*32 = 7.37
        rom[210] = 8'h08;    // exp(-1.438)*32 = 7.60 -> 8
        rom[211] = 8'h08;    // exp(-1.406)*32 = 7.84
        rom[212] = 8'h08;    // exp(-1.375)*32 = 8.09
        rom[213] = 8'h08;    // exp(-1.344)*32 = 8.35
        rom[214] = 8'h09;    // exp(-1.313)*32 = 8.62 -> 9
        rom[215] = 8'h09;    // exp(-1.281)*32 = 8.89
        rom[216] = 8'h09;    // exp(-1.250)*32 = 9.18
        rom[217] = 8'h09;    // exp(-1.219)*32 = 9.47
        rom[218] = 8'h0A;    // exp(-1.188)*32 = 9.77 -> 10
        rom[219] = 8'h0A;    // exp(-1.156)*32 = 10.08
        rom[220] = 8'h0A;    // exp(-1.125)*32 = 10.41
        rom[221] = 8'h0B;    // exp(-1.094)*32 = 10.74 -> 11
        rom[222] = 8'h0B;    // exp(-1.063)*32 = 11.08
        rom[223] = 8'h0B;    // exp(-1.031)*32 = 11.44
        rom[224] = 8'h0C;    // exp(-1.000)*32 = 11.77 -> 12
        rom[225] = 8'h0C;    // exp(-0.969)*32 = 12.15
        rom[226] = 8'h0D;    // exp(-0.938)*32 = 12.53 -> 13
        rom[227] = 8'h0D;    // exp(-0.906)*32 = 12.93
        rom[228] = 8'h0D;    // exp(-0.875)*32 = 13.34
        rom[229] = 8'h0E;    // exp(-0.844)*32 = 13.77 -> 14
        rom[230] = 8'h0E;    // exp(-0.813)*32 = 14.20
        rom[231] = 8'h0F;    // exp(-0.781)*32 = 14.66 -> 15
        rom[232] = 8'h0F;    // exp(-0.750)*32 = 15.12
        rom[233] = 8'h10;    // exp(-0.719)*32 = 15.60 -> 16
        rom[234] = 8'h10;    // exp(-0.688)*32 = 16.10
        rom[235] = 8'h11;    // exp(-0.656)*32 = 16.61 -> 17
        rom[236] = 8'h11;    // exp(-0.625)*32 = 17.14
        rom[237] = 8'h12;    // exp(-0.594)*32 = 17.69 -> 18
        rom[238] = 8'h12;    // exp(-0.563)*32 = 18.25
        rom[239] = 8'h13;    // exp(-0.531)*32 = 18.83 -> 19
        rom[240] = 8'h13;    // exp(-0.500)*32 = 19.41 -> 19
        rom[241] = 8'h14;    // exp(-0.469)*32 = 20.03 -> 20
        rom[242] = 8'h15;    // exp(-0.438)*32 = 20.66 -> 21
        rom[243] = 8'h15;    // exp(-0.406)*32 = 21.32
        rom[244] = 8'h16;    // exp(-0.375)*32 = 21.99 -> 22
        rom[245] = 8'h17;    // exp(-0.344)*32 = 22.69 -> 23
        rom[246] = 8'h17;    // exp(-0.313)*32 = 23.41
        rom[247] = 8'h18;    // exp(-0.281)*32 = 24.16 -> 24
        rom[248] = 8'h19;    // exp(-0.250)*32 = 24.92 -> 25
        rom[249] = 8'h1A;    // exp(-0.219)*32 = 25.71 -> 26
        rom[250] = 8'h1B;    // exp(-0.188)*32 = 26.54 -> 27
        rom[251] = 8'h1B;    // exp(-0.156)*32 = 27.39
        rom[252] = 8'h1C;    // exp(-0.125)*32 = 28.24 -> 28
        rom[253] = 8'h1D;    // exp(-0.094)*32 = 29.15 -> 29
        rom[254] = 8'h1E;    // exp(-0.063)*32 = 30.08 -> 30
        rom[255] = 8'h1F;    // exp(-0.031)*32 = 31.04 -> 31
    end

    // ----------------------------------------------------------------
    // Registered read (1-cycle latency)
    // ----------------------------------------------------------------
    always_ff @(posedge clk) begin
        data_out <= rom[addr];
    end

endmodule

`default_nettype wire
