// =============================================================================
// graph_sqrt_lut.sv - SQRT via 256-entry ROM lookup table
// Input:  x[7:0] signed int8
// Output: data_out[7:0] signed int8
// Formula: LUT[i] = clamp(round(sqrt(max(signed_i / 32, 0)) * 32), -128, 127)
// Scale: int8 maps to float via /32, so int8 range [-128,127] -> [-4.0, 3.97]
// Pipeline: 1-cycle registered output
// =============================================================================
`default_nettype none

module graph_sqrt_lut (
    input  wire        clk,
    input  wire  [7:0] addr,       // treated as signed int8 index
    output logic [7:0] data_out    // signed int8 SQRT result
);

    // 256-entry ROM - inferred as block RAM
    (* rom_style = "block" *)
    logic [7:0] rom [0:255];

    // ----------------------------------------------------------------
    // ROM initialization
    // LUT[i] = clamp(round(sqrt(max(signed_i/32.0, 0)) * 32.0), -128, 127)
    //
    // Key values (signed int8 index -> SQRT output):
    //   0   -> 0    (sqrt(0)*32 = 0)
    //   32  -> 32   (sqrt(1.0)*32 = 32)
    //   64  -> 45   (sqrt(2.0)*32 = 45.25)
    //  -128 -> 0    (negative input -> sqrt(0) = 0)
    // ----------------------------------------------------------------
    initial begin
        // Index 0 (signed 0): sqrt(0)*32 = 0
        rom[  0] = 8'h00;    // 0

        // Positive indices 1..127 (signed 1 to +127)
        // sqrt(n/32)*32 = 32*sqrt(n/32) = 5.6569*sqrt(n)
        rom[  1] = 8'h06;    // sqrt(0.031)*32 = 6
        rom[  2] = 8'h08;    // sqrt(0.063)*32 = 8
        rom[  3] = 8'h0A;    // sqrt(0.094)*32 = 10
        rom[  4] = 8'h0B;    // sqrt(0.125)*32 = 11
        rom[  5] = 8'h0D;    // sqrt(0.156)*32 = 13
        rom[  6] = 8'h0E;    // sqrt(0.188)*32 = 14
        rom[  7] = 8'h0F;    // sqrt(0.219)*32 = 15
        rom[  8] = 8'h10;    // sqrt(0.250)*32 = 16
        rom[  9] = 8'h11;    // sqrt(0.281)*32 = 17
        rom[ 10] = 8'h12;    // sqrt(0.313)*32 = 18
        rom[ 11] = 8'h13;    // sqrt(0.344)*32 = 19
        rom[ 12] = 8'h14;    // sqrt(0.375)*32 = 20
        rom[ 13] = 8'h14;    // sqrt(0.406)*32 = 20
        rom[ 14] = 8'h15;    // sqrt(0.438)*32 = 21
        rom[ 15] = 8'h16;    // sqrt(0.469)*32 = 22
        rom[ 16] = 8'h17;    // sqrt(0.500)*32 = 23
        rom[ 17] = 8'h17;    // sqrt(0.531)*32 = 23
        rom[ 18] = 8'h18;    // sqrt(0.563)*32 = 24
        rom[ 19] = 8'h19;    // sqrt(0.594)*32 = 25
        rom[ 20] = 8'h19;    // sqrt(0.625)*32 = 25
        rom[ 21] = 8'h1A;    // sqrt(0.656)*32 = 26
        rom[ 22] = 8'h1B;    // sqrt(0.688)*32 = 27
        rom[ 23] = 8'h1B;    // sqrt(0.719)*32 = 27
        rom[ 24] = 8'h1C;    // sqrt(0.750)*32 = 28
        rom[ 25] = 8'h1C;    // sqrt(0.781)*32 = 28
        rom[ 26] = 8'h1D;    // sqrt(0.813)*32 = 29
        rom[ 27] = 8'h1D;    // sqrt(0.844)*32 = 29
        rom[ 28] = 8'h1E;    // sqrt(0.875)*32 = 30
        rom[ 29] = 8'h1E;    // sqrt(0.906)*32 = 30
        rom[ 30] = 8'h1F;    // sqrt(0.938)*32 = 31
        rom[ 31] = 8'h1F;    // sqrt(0.969)*32 = 31
        rom[ 32] = 8'h20;    // sqrt(1.000)*32 = 32
        rom[ 33] = 8'h20;    // sqrt(1.031)*32 = 32
        rom[ 34] = 8'h21;    // sqrt(1.063)*32 = 33
        rom[ 35] = 8'h21;    // sqrt(1.094)*32 = 33
        rom[ 36] = 8'h22;    // sqrt(1.125)*32 = 34
        rom[ 37] = 8'h22;    // sqrt(1.156)*32 = 34
        rom[ 38] = 8'h23;    // sqrt(1.188)*32 = 35
        rom[ 39] = 8'h23;    // sqrt(1.219)*32 = 35
        rom[ 40] = 8'h24;    // sqrt(1.250)*32 = 36
        rom[ 41] = 8'h24;    // sqrt(1.281)*32 = 36
        rom[ 42] = 8'h25;    // sqrt(1.313)*32 = 37
        rom[ 43] = 8'h25;    // sqrt(1.344)*32 = 37
        rom[ 44] = 8'h26;    // sqrt(1.375)*32 = 38
        rom[ 45] = 8'h26;    // sqrt(1.406)*32 = 38
        rom[ 46] = 8'h26;    // sqrt(1.438)*32 = 38
        rom[ 47] = 8'h27;    // sqrt(1.469)*32 = 39
        rom[ 48] = 8'h27;    // sqrt(1.500)*32 = 39
        rom[ 49] = 8'h28;    // sqrt(1.531)*32 = 40
        rom[ 50] = 8'h28;    // sqrt(1.563)*32 = 40
        rom[ 51] = 8'h28;    // sqrt(1.594)*32 = 40
        rom[ 52] = 8'h29;    // sqrt(1.625)*32 = 41
        rom[ 53] = 8'h29;    // sqrt(1.656)*32 = 41
        rom[ 54] = 8'h2A;    // sqrt(1.688)*32 = 42
        rom[ 55] = 8'h2A;    // sqrt(1.719)*32 = 42
        rom[ 56] = 8'h2A;    // sqrt(1.750)*32 = 42
        rom[ 57] = 8'h2B;    // sqrt(1.781)*32 = 43
        rom[ 58] = 8'h2B;    // sqrt(1.813)*32 = 43
        rom[ 59] = 8'h2B;    // sqrt(1.844)*32 = 43
        rom[ 60] = 8'h2C;    // sqrt(1.875)*32 = 44
        rom[ 61] = 8'h2C;    // sqrt(1.906)*32 = 44
        rom[ 62] = 8'h2D;    // sqrt(1.938)*32 = 45
        rom[ 63] = 8'h2D;    // sqrt(1.969)*32 = 45
        rom[ 64] = 8'h2D;    // sqrt(2.000)*32 = 45
        rom[ 65] = 8'h2E;    // sqrt(2.031)*32 = 46
        rom[ 66] = 8'h2E;    // sqrt(2.063)*32 = 46
        rom[ 67] = 8'h2E;    // sqrt(2.094)*32 = 46
        rom[ 68] = 8'h2F;    // sqrt(2.125)*32 = 47
        rom[ 69] = 8'h2F;    // sqrt(2.156)*32 = 47
        rom[ 70] = 8'h2F;    // sqrt(2.188)*32 = 47
        rom[ 71] = 8'h30;    // sqrt(2.219)*32 = 48
        rom[ 72] = 8'h30;    // sqrt(2.250)*32 = 48
        rom[ 73] = 8'h30;    // sqrt(2.281)*32 = 48
        rom[ 74] = 8'h31;    // sqrt(2.313)*32 = 49
        rom[ 75] = 8'h31;    // sqrt(2.344)*32 = 49
        rom[ 76] = 8'h31;    // sqrt(2.375)*32 = 49
        rom[ 77] = 8'h32;    // sqrt(2.406)*32 = 50
        rom[ 78] = 8'h32;    // sqrt(2.438)*32 = 50
        rom[ 79] = 8'h32;    // sqrt(2.469)*32 = 50
        rom[ 80] = 8'h33;    // sqrt(2.500)*32 = 51
        rom[ 81] = 8'h33;    // sqrt(2.531)*32 = 51
        rom[ 82] = 8'h33;    // sqrt(2.563)*32 = 51
        rom[ 83] = 8'h34;    // sqrt(2.594)*32 = 52
        rom[ 84] = 8'h34;    // sqrt(2.625)*32 = 52
        rom[ 85] = 8'h34;    // sqrt(2.656)*32 = 52
        rom[ 86] = 8'h34;    // sqrt(2.688)*32 = 52
        rom[ 87] = 8'h35;    // sqrt(2.719)*32 = 53
        rom[ 88] = 8'h35;    // sqrt(2.750)*32 = 53
        rom[ 89] = 8'h35;    // sqrt(2.781)*32 = 53
        rom[ 90] = 8'h36;    // sqrt(2.813)*32 = 54
        rom[ 91] = 8'h36;    // sqrt(2.844)*32 = 54
        rom[ 92] = 8'h36;    // sqrt(2.875)*32 = 54
        rom[ 93] = 8'h37;    // sqrt(2.906)*32 = 55
        rom[ 94] = 8'h37;    // sqrt(2.938)*32 = 55
        rom[ 95] = 8'h37;    // sqrt(2.969)*32 = 55
        rom[ 96] = 8'h37;    // sqrt(3.000)*32 = 55
        rom[ 97] = 8'h38;    // sqrt(3.031)*32 = 56
        rom[ 98] = 8'h38;    // sqrt(3.063)*32 = 56
        rom[ 99] = 8'h38;    // sqrt(3.094)*32 = 56
        rom[100] = 8'h39;    // sqrt(3.125)*32 = 57
        rom[101] = 8'h39;    // sqrt(3.156)*32 = 57
        rom[102] = 8'h39;    // sqrt(3.188)*32 = 57
        rom[103] = 8'h39;    // sqrt(3.219)*32 = 57
        rom[104] = 8'h3A;    // sqrt(3.250)*32 = 58
        rom[105] = 8'h3A;    // sqrt(3.281)*32 = 58
        rom[106] = 8'h3A;    // sqrt(3.313)*32 = 58
        rom[107] = 8'h3B;    // sqrt(3.344)*32 = 59
        rom[108] = 8'h3B;    // sqrt(3.375)*32 = 59
        rom[109] = 8'h3B;    // sqrt(3.406)*32 = 59
        rom[110] = 8'h3B;    // sqrt(3.438)*32 = 59
        rom[111] = 8'h3C;    // sqrt(3.469)*32 = 60
        rom[112] = 8'h3C;    // sqrt(3.500)*32 = 60
        rom[113] = 8'h3C;    // sqrt(3.531)*32 = 60
        rom[114] = 8'h3C;    // sqrt(3.563)*32 = 60
        rom[115] = 8'h3D;    // sqrt(3.594)*32 = 61
        rom[116] = 8'h3D;    // sqrt(3.625)*32 = 61
        rom[117] = 8'h3D;    // sqrt(3.656)*32 = 61
        rom[118] = 8'h3D;    // sqrt(3.688)*32 = 61
        rom[119] = 8'h3E;    // sqrt(3.719)*32 = 62
        rom[120] = 8'h3E;    // sqrt(3.750)*32 = 62
        rom[121] = 8'h3E;    // sqrt(3.781)*32 = 62
        rom[122] = 8'h3E;    // sqrt(3.813)*32 = 62
        rom[123] = 8'h3F;    // sqrt(3.844)*32 = 63
        rom[124] = 8'h3F;    // sqrt(3.875)*32 = 63
        rom[125] = 8'h3F;    // sqrt(3.906)*32 = 63
        rom[126] = 8'h3F;    // sqrt(3.938)*32 = 63
        rom[127] = 8'h40;    // sqrt(3.969)*32 = 64

        // Negative indices 128..255 (signed -128 to -1)
        // All negative inputs: max(signed_i/32, 0) = 0
        // sqrt(0)*32 = 0
        rom[128] = 8'h00;
        rom[129] = 8'h00;
        rom[130] = 8'h00;
        rom[131] = 8'h00;
        rom[132] = 8'h00;
        rom[133] = 8'h00;
        rom[134] = 8'h00;
        rom[135] = 8'h00;
        rom[136] = 8'h00;
        rom[137] = 8'h00;
        rom[138] = 8'h00;
        rom[139] = 8'h00;
        rom[140] = 8'h00;
        rom[141] = 8'h00;
        rom[142] = 8'h00;
        rom[143] = 8'h00;
        rom[144] = 8'h00;
        rom[145] = 8'h00;
        rom[146] = 8'h00;
        rom[147] = 8'h00;
        rom[148] = 8'h00;
        rom[149] = 8'h00;
        rom[150] = 8'h00;
        rom[151] = 8'h00;
        rom[152] = 8'h00;
        rom[153] = 8'h00;
        rom[154] = 8'h00;
        rom[155] = 8'h00;
        rom[156] = 8'h00;
        rom[157] = 8'h00;
        rom[158] = 8'h00;
        rom[159] = 8'h00;
        rom[160] = 8'h00;
        rom[161] = 8'h00;
        rom[162] = 8'h00;
        rom[163] = 8'h00;
        rom[164] = 8'h00;
        rom[165] = 8'h00;
        rom[166] = 8'h00;
        rom[167] = 8'h00;
        rom[168] = 8'h00;
        rom[169] = 8'h00;
        rom[170] = 8'h00;
        rom[171] = 8'h00;
        rom[172] = 8'h00;
        rom[173] = 8'h00;
        rom[174] = 8'h00;
        rom[175] = 8'h00;
        rom[176] = 8'h00;
        rom[177] = 8'h00;
        rom[178] = 8'h00;
        rom[179] = 8'h00;
        rom[180] = 8'h00;
        rom[181] = 8'h00;
        rom[182] = 8'h00;
        rom[183] = 8'h00;
        rom[184] = 8'h00;
        rom[185] = 8'h00;
        rom[186] = 8'h00;
        rom[187] = 8'h00;
        rom[188] = 8'h00;
        rom[189] = 8'h00;
        rom[190] = 8'h00;
        rom[191] = 8'h00;
        rom[192] = 8'h00;
        rom[193] = 8'h00;
        rom[194] = 8'h00;
        rom[195] = 8'h00;
        rom[196] = 8'h00;
        rom[197] = 8'h00;
        rom[198] = 8'h00;
        rom[199] = 8'h00;
        rom[200] = 8'h00;
        rom[201] = 8'h00;
        rom[202] = 8'h00;
        rom[203] = 8'h00;
        rom[204] = 8'h00;
        rom[205] = 8'h00;
        rom[206] = 8'h00;
        rom[207] = 8'h00;
        rom[208] = 8'h00;
        rom[209] = 8'h00;
        rom[210] = 8'h00;
        rom[211] = 8'h00;
        rom[212] = 8'h00;
        rom[213] = 8'h00;
        rom[214] = 8'h00;
        rom[215] = 8'h00;
        rom[216] = 8'h00;
        rom[217] = 8'h00;
        rom[218] = 8'h00;
        rom[219] = 8'h00;
        rom[220] = 8'h00;
        rom[221] = 8'h00;
        rom[222] = 8'h00;
        rom[223] = 8'h00;
        rom[224] = 8'h00;
        rom[225] = 8'h00;
        rom[226] = 8'h00;
        rom[227] = 8'h00;
        rom[228] = 8'h00;
        rom[229] = 8'h00;
        rom[230] = 8'h00;
        rom[231] = 8'h00;
        rom[232] = 8'h00;
        rom[233] = 8'h00;
        rom[234] = 8'h00;
        rom[235] = 8'h00;
        rom[236] = 8'h00;
        rom[237] = 8'h00;
        rom[238] = 8'h00;
        rom[239] = 8'h00;
        rom[240] = 8'h00;
        rom[241] = 8'h00;
        rom[242] = 8'h00;
        rom[243] = 8'h00;
        rom[244] = 8'h00;
        rom[245] = 8'h00;
        rom[246] = 8'h00;
        rom[247] = 8'h00;
        rom[248] = 8'h00;
        rom[249] = 8'h00;
        rom[250] = 8'h00;
        rom[251] = 8'h00;
        rom[252] = 8'h00;
        rom[253] = 8'h00;
        rom[254] = 8'h00;
        rom[255] = 8'h00;
    end

    // ----------------------------------------------------------------
    // Registered read (1-cycle latency)
    // ----------------------------------------------------------------
    always_ff @(posedge clk) begin
        data_out <= rom[addr];
    end

endmodule

`default_nettype wire
