// =============================================================================
// graph_log_lut.sv - LOG (natural log) via 256-entry ROM lookup table
// Input:  x[7:0] signed int8
// Output: data_out[7:0] signed int8
// Formula: LUT[i] = clamp(round(log(max(signed_i / 32, 0.001)) * 32), -128, 127)
// Scale: int8 maps to float via /32, so int8 range [-128,127] -> [-4.0, 3.97]
// Pipeline: 1-cycle registered output
// =============================================================================
`default_nettype none

module graph_log_lut (
    input  wire        clk,
    input  wire  [7:0] addr,       // treated as signed int8 index
    output logic [7:0] data_out    // signed int8 LOG result
);

    // 256-entry ROM - inferred as block RAM
    (* rom_style = "block" *)
    logic [7:0] rom [0:255];

    // ----------------------------------------------------------------
    // ROM initialization
    // LUT[i] = clamp(round(log(max(signed_i/32.0, 0.001)) * 32.0), -128, 127)
    //
    // Key values (signed int8 index -> LOG output):
    //   0   -> -128 (log(0.001)*32 = -221 -> clamped)
    //   32  -> 0    (log(1.0)*32 = 0)
    //   64  -> 22   (log(2.0)*32 = 22.18)
    //  -128 -> -128 (negative input -> log(0.001) -> clamped)
    // ----------------------------------------------------------------
    initial begin
        // Index 0 (signed 0): max(0/32, 0.001)=0.001, log(0.001)*32=-221 -> -128
        rom[  0] = 8'h80;    // -128

        // Positive indices 1..127 (signed 1 to +127)
        // x_float = i/32.0, range [0.03125, 3.97]
        rom[  1] = 8'h91;    // log(0.031)*32 = -111
        rom[  2] = 8'hA7;    // log(0.063)*32 = -89
        rom[  3] = 8'hB4;    // log(0.094)*32 = -76
        rom[  4] = 8'hBD;    // log(0.125)*32 = -67
        rom[  5] = 8'hC5;    // log(0.156)*32 = -59
        rom[  6] = 8'hCA;    // log(0.188)*32 = -54
        rom[  7] = 8'hCF;    // log(0.219)*32 = -49
        rom[  8] = 8'hD4;    // log(0.250)*32 = -44
        rom[  9] = 8'hD7;    // log(0.281)*32 = -41
        rom[ 10] = 8'hDB;    // log(0.313)*32 = -37
        rom[ 11] = 8'hDE;    // log(0.344)*32 = -34
        rom[ 12] = 8'hE1;    // log(0.375)*32 = -31
        rom[ 13] = 8'hE3;    // log(0.406)*32 = -29
        rom[ 14] = 8'hE6;    // log(0.438)*32 = -26
        rom[ 15] = 8'hE8;    // log(0.469)*32 = -24
        rom[ 16] = 8'hEA;    // log(0.500)*32 = -22
        rom[ 17] = 8'hEC;    // log(0.531)*32 = -20
        rom[ 18] = 8'hEE;    // log(0.563)*32 = -18
        rom[ 19] = 8'hEF;    // log(0.594)*32 = -17
        rom[ 20] = 8'hF1;    // log(0.625)*32 = -15
        rom[ 21] = 8'hF3;    // log(0.656)*32 = -13
        rom[ 22] = 8'hF4;    // log(0.688)*32 = -12
        rom[ 23] = 8'hF5;    // log(0.719)*32 = -11
        rom[ 24] = 8'hF7;    // log(0.750)*32 = -9
        rom[ 25] = 8'hF8;    // log(0.781)*32 = -8
        rom[ 26] = 8'hF9;    // log(0.813)*32 = -7
        rom[ 27] = 8'hFB;    // log(0.844)*32 = -5
        rom[ 28] = 8'hFC;    // log(0.875)*32 = -4
        rom[ 29] = 8'hFD;    // log(0.906)*32 = -3
        rom[ 30] = 8'hFE;    // log(0.938)*32 = -2
        rom[ 31] = 8'hFF;    // log(0.969)*32 = -1
        rom[ 32] = 8'h00;    // log(1.000)*32 = 0
        rom[ 33] = 8'h01;    // log(1.031)*32 = 1
        rom[ 34] = 8'h02;    // log(1.063)*32 = 2
        rom[ 35] = 8'h03;    // log(1.094)*32 = 3
        rom[ 36] = 8'h04;    // log(1.125)*32 = 4
        rom[ 37] = 8'h05;    // log(1.156)*32 = 5
        rom[ 38] = 8'h05;    // log(1.188)*32 = 5
        rom[ 39] = 8'h06;    // log(1.219)*32 = 6
        rom[ 40] = 8'h07;    // log(1.250)*32 = 7
        rom[ 41] = 8'h08;    // log(1.281)*32 = 8
        rom[ 42] = 8'h09;    // log(1.313)*32 = 9
        rom[ 43] = 8'h09;    // log(1.344)*32 = 9
        rom[ 44] = 8'h0A;    // log(1.375)*32 = 10
        rom[ 45] = 8'h0B;    // log(1.406)*32 = 11
        rom[ 46] = 8'h0C;    // log(1.438)*32 = 12
        rom[ 47] = 8'h0C;    // log(1.469)*32 = 12
        rom[ 48] = 8'h0D;    // log(1.500)*32 = 13
        rom[ 49] = 8'h0E;    // log(1.531)*32 = 14
        rom[ 50] = 8'h0E;    // log(1.563)*32 = 14
        rom[ 51] = 8'h0F;    // log(1.594)*32 = 15
        rom[ 52] = 8'h10;    // log(1.625)*32 = 16
        rom[ 53] = 8'h10;    // log(1.656)*32 = 16
        rom[ 54] = 8'h11;    // log(1.688)*32 = 17
        rom[ 55] = 8'h11;    // log(1.719)*32 = 17
        rom[ 56] = 8'h12;    // log(1.750)*32 = 18
        rom[ 57] = 8'h12;    // log(1.781)*32 = 18
        rom[ 58] = 8'h13;    // log(1.813)*32 = 19
        rom[ 59] = 8'h14;    // log(1.844)*32 = 20
        rom[ 60] = 8'h14;    // log(1.875)*32 = 20
        rom[ 61] = 8'h15;    // log(1.906)*32 = 21
        rom[ 62] = 8'h15;    // log(1.938)*32 = 21
        rom[ 63] = 8'h16;    // log(1.969)*32 = 22
        rom[ 64] = 8'h16;    // log(2.000)*32 = 22
        rom[ 65] = 8'h17;    // log(2.031)*32 = 23
        rom[ 66] = 8'h17;    // log(2.063)*32 = 23
        rom[ 67] = 8'h18;    // log(2.094)*32 = 24
        rom[ 68] = 8'h18;    // log(2.125)*32 = 24
        rom[ 69] = 8'h19;    // log(2.156)*32 = 25
        rom[ 70] = 8'h19;    // log(2.188)*32 = 25
        rom[ 71] = 8'h19;    // log(2.219)*32 = 25
        rom[ 72] = 8'h1A;    // log(2.250)*32 = 26
        rom[ 73] = 8'h1A;    // log(2.281)*32 = 26
        rom[ 74] = 8'h1B;    // log(2.313)*32 = 27
        rom[ 75] = 8'h1B;    // log(2.344)*32 = 27
        rom[ 76] = 8'h1C;    // log(2.375)*32 = 28
        rom[ 77] = 8'h1C;    // log(2.406)*32 = 28
        rom[ 78] = 8'h1D;    // log(2.438)*32 = 29
        rom[ 79] = 8'h1D;    // log(2.469)*32 = 29
        rom[ 80] = 8'h1D;    // log(2.500)*32 = 29
        rom[ 81] = 8'h1E;    // log(2.531)*32 = 30
        rom[ 82] = 8'h1E;    // log(2.563)*32 = 30
        rom[ 83] = 8'h1E;    // log(2.594)*32 = 30
        rom[ 84] = 8'h1F;    // log(2.625)*32 = 31
        rom[ 85] = 8'h1F;    // log(2.656)*32 = 31
        rom[ 86] = 8'h20;    // log(2.688)*32 = 32
        rom[ 87] = 8'h20;    // log(2.719)*32 = 32
        rom[ 88] = 8'h20;    // log(2.750)*32 = 32
        rom[ 89] = 8'h21;    // log(2.781)*32 = 33
        rom[ 90] = 8'h21;    // log(2.813)*32 = 33
        rom[ 91] = 8'h21;    // log(2.844)*32 = 33
        rom[ 92] = 8'h22;    // log(2.875)*32 = 34
        rom[ 93] = 8'h22;    // log(2.906)*32 = 34
        rom[ 94] = 8'h22;    // log(2.938)*32 = 34
        rom[ 95] = 8'h23;    // log(2.969)*32 = 35
        rom[ 96] = 8'h23;    // log(3.000)*32 = 35
        rom[ 97] = 8'h23;    // log(3.031)*32 = 35
        rom[ 98] = 8'h24;    // log(3.063)*32 = 36
        rom[ 99] = 8'h24;    // log(3.094)*32 = 36
        rom[100] = 8'h24;    // log(3.125)*32 = 36
        rom[101] = 8'h25;    // log(3.156)*32 = 37
        rom[102] = 8'h25;    // log(3.188)*32 = 37
        rom[103] = 8'h25;    // log(3.219)*32 = 37
        rom[104] = 8'h26;    // log(3.250)*32 = 38
        rom[105] = 8'h26;    // log(3.281)*32 = 38
        rom[106] = 8'h26;    // log(3.313)*32 = 38
        rom[107] = 8'h27;    // log(3.344)*32 = 39
        rom[108] = 8'h27;    // log(3.375)*32 = 39
        rom[109] = 8'h27;    // log(3.406)*32 = 39
        rom[110] = 8'h28;    // log(3.438)*32 = 40
        rom[111] = 8'h28;    // log(3.469)*32 = 40
        rom[112] = 8'h28;    // log(3.500)*32 = 40
        rom[113] = 8'h28;    // log(3.531)*32 = 40
        rom[114] = 8'h29;    // log(3.563)*32 = 41
        rom[115] = 8'h29;    // log(3.594)*32 = 41
        rom[116] = 8'h29;    // log(3.625)*32 = 41
        rom[117] = 8'h29;    // log(3.656)*32 = 41
        rom[118] = 8'h2A;    // log(3.688)*32 = 42
        rom[119] = 8'h2A;    // log(3.719)*32 = 42
        rom[120] = 8'h2A;    // log(3.750)*32 = 42
        rom[121] = 8'h2B;    // log(3.781)*32 = 43
        rom[122] = 8'h2B;    // log(3.813)*32 = 43
        rom[123] = 8'h2B;    // log(3.844)*32 = 43
        rom[124] = 8'h2B;    // log(3.875)*32 = 43
        rom[125] = 8'h2C;    // log(3.906)*32 = 44
        rom[126] = 8'h2C;    // log(3.938)*32 = 44
        rom[127] = 8'h2C;    // log(3.969)*32 = 44

        // Negative indices 128..255 (signed -128 to -1)
        // All negative inputs: max(signed_i/32, 0.001) = 0.001
        // log(0.001)*32 = -221.05 -> clamped to -128
        rom[128] = 8'h80;    // -128
        rom[129] = 8'h80;
        rom[130] = 8'h80;
        rom[131] = 8'h80;
        rom[132] = 8'h80;
        rom[133] = 8'h80;
        rom[134] = 8'h80;
        rom[135] = 8'h80;
        rom[136] = 8'h80;
        rom[137] = 8'h80;
        rom[138] = 8'h80;
        rom[139] = 8'h80;
        rom[140] = 8'h80;
        rom[141] = 8'h80;
        rom[142] = 8'h80;
        rom[143] = 8'h80;
        rom[144] = 8'h80;
        rom[145] = 8'h80;
        rom[146] = 8'h80;
        rom[147] = 8'h80;
        rom[148] = 8'h80;
        rom[149] = 8'h80;
        rom[150] = 8'h80;
        rom[151] = 8'h80;
        rom[152] = 8'h80;
        rom[153] = 8'h80;
        rom[154] = 8'h80;
        rom[155] = 8'h80;
        rom[156] = 8'h80;
        rom[157] = 8'h80;
        rom[158] = 8'h80;
        rom[159] = 8'h80;
        rom[160] = 8'h80;
        rom[161] = 8'h80;
        rom[162] = 8'h80;
        rom[163] = 8'h80;
        rom[164] = 8'h80;
        rom[165] = 8'h80;
        rom[166] = 8'h80;
        rom[167] = 8'h80;
        rom[168] = 8'h80;
        rom[169] = 8'h80;
        rom[170] = 8'h80;
        rom[171] = 8'h80;
        rom[172] = 8'h80;
        rom[173] = 8'h80;
        rom[174] = 8'h80;
        rom[175] = 8'h80;
        rom[176] = 8'h80;
        rom[177] = 8'h80;
        rom[178] = 8'h80;
        rom[179] = 8'h80;
        rom[180] = 8'h80;
        rom[181] = 8'h80;
        rom[182] = 8'h80;
        rom[183] = 8'h80;
        rom[184] = 8'h80;
        rom[185] = 8'h80;
        rom[186] = 8'h80;
        rom[187] = 8'h80;
        rom[188] = 8'h80;
        rom[189] = 8'h80;
        rom[190] = 8'h80;
        rom[191] = 8'h80;
        rom[192] = 8'h80;
        rom[193] = 8'h80;
        rom[194] = 8'h80;
        rom[195] = 8'h80;
        rom[196] = 8'h80;
        rom[197] = 8'h80;
        rom[198] = 8'h80;
        rom[199] = 8'h80;
        rom[200] = 8'h80;
        rom[201] = 8'h80;
        rom[202] = 8'h80;
        rom[203] = 8'h80;
        rom[204] = 8'h80;
        rom[205] = 8'h80;
        rom[206] = 8'h80;
        rom[207] = 8'h80;
        rom[208] = 8'h80;
        rom[209] = 8'h80;
        rom[210] = 8'h80;
        rom[211] = 8'h80;
        rom[212] = 8'h80;
        rom[213] = 8'h80;
        rom[214] = 8'h80;
        rom[215] = 8'h80;
        rom[216] = 8'h80;
        rom[217] = 8'h80;
        rom[218] = 8'h80;
        rom[219] = 8'h80;
        rom[220] = 8'h80;
        rom[221] = 8'h80;
        rom[222] = 8'h80;
        rom[223] = 8'h80;
        rom[224] = 8'h80;
        rom[225] = 8'h80;
        rom[226] = 8'h80;
        rom[227] = 8'h80;
        rom[228] = 8'h80;
        rom[229] = 8'h80;
        rom[230] = 8'h80;
        rom[231] = 8'h80;
        rom[232] = 8'h80;
        rom[233] = 8'h80;
        rom[234] = 8'h80;
        rom[235] = 8'h80;
        rom[236] = 8'h80;
        rom[237] = 8'h80;
        rom[238] = 8'h80;
        rom[239] = 8'h80;
        rom[240] = 8'h80;
        rom[241] = 8'h80;
        rom[242] = 8'h80;
        rom[243] = 8'h80;
        rom[244] = 8'h80;
        rom[245] = 8'h80;
        rom[246] = 8'h80;
        rom[247] = 8'h80;
        rom[248] = 8'h80;
        rom[249] = 8'h80;
        rom[250] = 8'h80;
        rom[251] = 8'h80;
        rom[252] = 8'h80;
        rom[253] = 8'h80;
        rom[254] = 8'h80;
        rom[255] = 8'h80;
    end

    // ----------------------------------------------------------------
    // Registered read (1-cycle latency)
    // ----------------------------------------------------------------
    always_ff @(posedge clk) begin
        data_out <= rom[addr];
    end

endmodule

`default_nettype wire
