// =============================================================================
// recip_lut.sv - Reciprocal (1/x) approximation via 256-entry ROM
// Input:  x[15:0] unsigned (sum from reduce_sum, Q8.8 format)
// Output: recip_out[15:0] unsigned (Q0.16 format, so 1/256 maps to 256)
// Index:  top 8 bits of x are used as LUT index
// LUT:    recip_lut[i] = round(65536 / max(i, 1)) with i=0 special-cased
// Includes optional Newton-Raphson refinement for better accuracy
// Pipeline: 1-cycle registered (LUT only), or 2-cycle with NR refinement
// =============================================================================
import npu_pkg::*;
import fixed_pkg::*;

module recip_lut (
    input  logic        clk,
    input  logic [7:0]  addr,       // top 8 bits of the 16-bit sum
    output logic [15:0] data_out    // Q0.16 reciprocal
);

    // 256-entry ROM - inferred as block RAM
    (* rom_style = "block" *)
    logic [15:0] rom [0:255];

    // ----------------------------------------------------------------
    // ROM initialization
    // recip_lut[i] = round(65536 / max(i, 1))
    // i=0 -> special case: max value (65535)
    // i=1 -> 65536/1 = 65536 -> clamped to 65535
    // i=2 -> 65536/2 = 32768
    // i=128 -> 65536/128 = 512
    // i=255 -> 65536/255 = 257
    // ----------------------------------------------------------------
    initial begin
        rom[  0] = 16'hFFFF;  // special: 1/0 = max
        rom[  1] = 16'hFFFF;  // 65536/1 clamped
        rom[  2] = 16'd32768; // 65536/2
        rom[  3] = 16'd21845;
        rom[  4] = 16'd16384;
        rom[  5] = 16'd13107;
        rom[  6] = 16'd10923;
        rom[  7] = 16'd9362;
        rom[  8] = 16'd8192;
        rom[  9] = 16'd7282;
        rom[ 10] = 16'd6554;
        rom[ 11] = 16'd5958;
        rom[ 12] = 16'd5461;
        rom[ 13] = 16'd5041;
        rom[ 14] = 16'd4681;
        rom[ 15] = 16'd4369;
        rom[ 16] = 16'd4096;
        rom[ 17] = 16'd3855;
        rom[ 18] = 16'd3641;
        rom[ 19] = 16'd3449;
        rom[ 20] = 16'd3277;
        rom[ 21] = 16'd3121;
        rom[ 22] = 16'd2979;
        rom[ 23] = 16'd2849;
        rom[ 24] = 16'd2731;
        rom[ 25] = 16'd2621;
        rom[ 26] = 16'd2521;
        rom[ 27] = 16'd2427;
        rom[ 28] = 16'd2341;
        rom[ 29] = 16'd2260;
        rom[ 30] = 16'd2185;
        rom[ 31] = 16'd2114;
        rom[ 32] = 16'd2048;
        rom[ 33] = 16'd1986;
        rom[ 34] = 16'd1928;
        rom[ 35] = 16'd1872;
        rom[ 36] = 16'd1820;
        rom[ 37] = 16'd1771;
        rom[ 38] = 16'd1725;
        rom[ 39] = 16'd1680;
        rom[ 40] = 16'd1638;
        rom[ 41] = 16'd1598;
        rom[ 42] = 16'd1560;
        rom[ 43] = 16'd1524;
        rom[ 44] = 16'd1489;
        rom[ 45] = 16'd1456;
        rom[ 46] = 16'd1425;
        rom[ 47] = 16'd1394;
        rom[ 48] = 16'd1365;
        rom[ 49] = 16'd1337;
        rom[ 50] = 16'd1311;
        rom[ 51] = 16'd1285;
        rom[ 52] = 16'd1260;
        rom[ 53] = 16'd1237;
        rom[ 54] = 16'd1214;
        rom[ 55] = 16'd1192;
        rom[ 56] = 16'd1170;
        rom[ 57] = 16'd1150;
        rom[ 58] = 16'd1130;
        rom[ 59] = 16'd1111;
        rom[ 60] = 16'd1092;
        rom[ 61] = 16'd1074;
        rom[ 62] = 16'd1057;
        rom[ 63] = 16'd1040;
        rom[ 64] = 16'd1024;
        rom[ 65] = 16'd1008;
        rom[ 66] = 16'd993;
        rom[ 67] = 16'd978;
        rom[ 68] = 16'd964;
        rom[ 69] = 16'd950;
        rom[ 70] = 16'd936;
        rom[ 71] = 16'd923;
        rom[ 72] = 16'd910;
        rom[ 73] = 16'd898;
        rom[ 74] = 16'd886;
        rom[ 75] = 16'd874;
        rom[ 76] = 16'd862;
        rom[ 77] = 16'd851;
        rom[ 78] = 16'd840;
        rom[ 79] = 16'd830;
        rom[ 80] = 16'd819;
        rom[ 81] = 16'd809;
        rom[ 82] = 16'd799;
        rom[ 83] = 16'd789;
        rom[ 84] = 16'd780;
        rom[ 85] = 16'd771;
        rom[ 86] = 16'd762;
        rom[ 87] = 16'd753;
        rom[ 88] = 16'd745;
        rom[ 89] = 16'd736;
        rom[ 90] = 16'd728;
        rom[ 91] = 16'd720;
        rom[ 92] = 16'd712;
        rom[ 93] = 16'd705;
        rom[ 94] = 16'd697;
        rom[ 95] = 16'd690;
        rom[ 96] = 16'd683;
        rom[ 97] = 16'd676;
        rom[ 98] = 16'd669;
        rom[ 99] = 16'd662;
        rom[100] = 16'd655;
        rom[101] = 16'd649;
        rom[102] = 16'd643;
        rom[103] = 16'd636;
        rom[104] = 16'd630;
        rom[105] = 16'd624;
        rom[106] = 16'd618;
        rom[107] = 16'd612;
        rom[108] = 16'd607;
        rom[109] = 16'd601;
        rom[110] = 16'd596;
        rom[111] = 16'd591;
        rom[112] = 16'd585;
        rom[113] = 16'd580;
        rom[114] = 16'd575;
        rom[115] = 16'd570;
        rom[116] = 16'd565;
        rom[117] = 16'd560;
        rom[118] = 16'd555;
        rom[119] = 16'd551;
        rom[120] = 16'd546;
        rom[121] = 16'd542;
        rom[122] = 16'd537;
        rom[123] = 16'd533;
        rom[124] = 16'd529;
        rom[125] = 16'd524;
        rom[126] = 16'd520;
        rom[127] = 16'd516;
        rom[128] = 16'd512;
        rom[129] = 16'd508;
        rom[130] = 16'd504;
        rom[131] = 16'd500;
        rom[132] = 16'd497;
        rom[133] = 16'd493;
        rom[134] = 16'd489;
        rom[135] = 16'd486;
        rom[136] = 16'd482;
        rom[137] = 16'd479;
        rom[138] = 16'd475;
        rom[139] = 16'd472;
        rom[140] = 16'd468;
        rom[141] = 16'd465;
        rom[142] = 16'd462;
        rom[143] = 16'd458;
        rom[144] = 16'd455;
        rom[145] = 16'd452;
        rom[146] = 16'd449;
        rom[147] = 16'd446;
        rom[148] = 16'd443;
        rom[149] = 16'd440;
        rom[150] = 16'd437;
        rom[151] = 16'd434;
        rom[152] = 16'd431;
        rom[153] = 16'd428;
        rom[154] = 16'd426;
        rom[155] = 16'd423;
        rom[156] = 16'd420;
        rom[157] = 16'd418;
        rom[158] = 16'd415;
        rom[159] = 16'd412;
        rom[160] = 16'd410;
        rom[161] = 16'd407;
        rom[162] = 16'd405;
        rom[163] = 16'd402;
        rom[164] = 16'd400;
        rom[165] = 16'd397;
        rom[166] = 16'd395;
        rom[167] = 16'd393;
        rom[168] = 16'd390;
        rom[169] = 16'd388;
        rom[170] = 16'd386;
        rom[171] = 16'd383;
        rom[172] = 16'd381;
        rom[173] = 16'd379;
        rom[174] = 16'd377;
        rom[175] = 16'd375;
        rom[176] = 16'd372;
        rom[177] = 16'd370;
        rom[178] = 16'd368;
        rom[179] = 16'd366;
        rom[180] = 16'd364;
        rom[181] = 16'd362;
        rom[182] = 16'd360;
        rom[183] = 16'd358;
        rom[184] = 16'd356;
        rom[185] = 16'd354;
        rom[186] = 16'd352;
        rom[187] = 16'd351;
        rom[188] = 16'd349;
        rom[189] = 16'd347;
        rom[190] = 16'd345;
        rom[191] = 16'd343;
        rom[192] = 16'd341;
        rom[193] = 16'd340;
        rom[194] = 16'd338;
        rom[195] = 16'd336;
        rom[196] = 16'd334;
        rom[197] = 16'd333;
        rom[198] = 16'd331;
        rom[199] = 16'd329;
        rom[200] = 16'd328;
        rom[201] = 16'd326;
        rom[202] = 16'd325;
        rom[203] = 16'd323;
        rom[204] = 16'd321;
        rom[205] = 16'd320;
        rom[206] = 16'd318;
        rom[207] = 16'd317;
        rom[208] = 16'd315;
        rom[209] = 16'd314;
        rom[210] = 16'd312;
        rom[211] = 16'd311;
        rom[212] = 16'd309;
        rom[213] = 16'd308;
        rom[214] = 16'd306;
        rom[215] = 16'd305;
        rom[216] = 16'd303;
        rom[217] = 16'd302;
        rom[218] = 16'd301;
        rom[219] = 16'd299;
        rom[220] = 16'd298;
        rom[221] = 16'd297;
        rom[222] = 16'd295;
        rom[223] = 16'd294;
        rom[224] = 16'd293;
        rom[225] = 16'd291;
        rom[226] = 16'd290;
        rom[227] = 16'd289;
        rom[228] = 16'd288;
        rom[229] = 16'd286;
        rom[230] = 16'd285;
        rom[231] = 16'd284;
        rom[232] = 16'd282;
        rom[233] = 16'd281;
        rom[234] = 16'd280;
        rom[235] = 16'd279;
        rom[236] = 16'd278;
        rom[237] = 16'd276;
        rom[238] = 16'd275;
        rom[239] = 16'd274;
        rom[240] = 16'd273;
        rom[241] = 16'd272;
        rom[242] = 16'd271;
        rom[243] = 16'd270;
        rom[244] = 16'd269;
        rom[245] = 16'd267;
        rom[246] = 16'd266;
        rom[247] = 16'd265;
        rom[248] = 16'd264;
        rom[249] = 16'd263;
        rom[250] = 16'd262;
        rom[251] = 16'd261;
        rom[252] = 16'd260;
        rom[253] = 16'd259;
        rom[254] = 16'd258;
        rom[255] = 16'd257;
    end

    // ----------------------------------------------------------------
    // Registered read (1-cycle latency)
    // ----------------------------------------------------------------
    always_ff @(posedge clk) begin
        data_out <= rom[addr];
    end

endmodule
