// =============================================================================
// exp_lut.sv - Exponential approximation via 256-entry ROM lookup table
// Input:  x[7:0] signed (representing x - max, so always <= 0 in [-128, 0])
// Output: exp_out[15:0] unsigned Q8.8 fixed-point
//         exp(0) = 256, exp(-1) ~ 248, exp(-128) ~ 0
// LUT: exp_out[i] = clamp(round(256 * exp(signed(i) / 32.0)), 0, 65535)
// Pipeline: 1-cycle registered output
// =============================================================================
import npu_pkg::*;
import fixed_pkg::*;

module exp_lut (
    input  logic        clk,
    input  logic [7:0]  addr,       // treated as signed index for the function
    output logic [15:0] data_out    // Q8.8 unsigned result
);

    // 256-entry ROM - inferred as block RAM
    (* rom_style = "block" *)
    logic [15:0] rom [0:255];

    // ----------------------------------------------------------------
    // ROM initialization
    // Values: exp_out[i] = clamp(round(256 * exp(signed_i / 32.0)), 0, 65535)
    // where signed_i = (i < 128) ? i : i - 256
    // For softmax: input is (x - max), so signed_i <= 0 for valid inputs
    //   signed_i =   0 -> exp(0)    = 256
    //   signed_i =  -1 -> exp(-1/32)= 248
    //   signed_i = -32 -> exp(-1)   = 94
    //   signed_i = -128-> exp(-4)   = 5
    // Placeholder values - regenerate with make_lut.py for full precision
    // ----------------------------------------------------------------
    initial begin
        // Positive side (signed 0..127): exp(i/32)*256, clamped to 16-bit
        rom[  0] = 16'd256;    // exp(0/32)*256 = 256
        rom[  1] = 16'd264;    // exp(1/32)*256
        rom[  2] = 16'd272;    // exp(2/32)*256
        rom[  3] = 16'd281;
        rom[  4] = 16'd289;
        rom[  5] = 16'd298;
        rom[  6] = 16'd308;
        rom[  7] = 16'd317;
        rom[  8] = 16'd327;    // exp(0.25)*256 = 329
        rom[  9] = 16'd337;
        rom[ 10] = 16'd348;
        rom[ 11] = 16'd358;
        rom[ 12] = 16'd369;
        rom[ 13] = 16'd381;
        rom[ 14] = 16'd392;
        rom[ 15] = 16'd404;
        rom[ 16] = 16'd417;    // exp(0.5)*256 = 422
        rom[ 17] = 16'd430;
        rom[ 18] = 16'd443;
        rom[ 19] = 16'd456;
        rom[ 20] = 16'd470;
        rom[ 21] = 16'd485;
        rom[ 22] = 16'd500;
        rom[ 23] = 16'd515;
        rom[ 24] = 16'd531;    // exp(0.75)*256 = 542
        rom[ 25] = 16'd548;
        rom[ 26] = 16'd565;
        rom[ 27] = 16'd582;
        rom[ 28] = 16'd600;
        rom[ 29] = 16'd618;
        rom[ 30] = 16'd637;
        rom[ 31] = 16'd657;
        rom[ 32] = 16'd696;    // exp(1.0)*256 = 696
        rom[ 33] = 16'd718;
        rom[ 34] = 16'd740;
        rom[ 35] = 16'd763;
        rom[ 36] = 16'd786;
        rom[ 37] = 16'd810;
        rom[ 38] = 16'd835;
        rom[ 39] = 16'd861;
        rom[ 40] = 16'd887;
        rom[ 41] = 16'd914;
        rom[ 42] = 16'd942;
        rom[ 43] = 16'd971;
        rom[ 44] = 16'd1001;
        rom[ 45] = 16'd1032;
        rom[ 46] = 16'd1063;
        rom[ 47] = 16'd1096;
        rom[ 48] = 16'd1130;   // exp(1.5)*256 = 1147
        rom[ 49] = 16'd1164;
        rom[ 50] = 16'd1200;
        rom[ 51] = 16'd1237;
        rom[ 52] = 16'd1275;
        rom[ 53] = 16'd1314;
        rom[ 54] = 16'd1354;
        rom[ 55] = 16'd1396;
        rom[ 56] = 16'd1438;
        rom[ 57] = 16'd1482;
        rom[ 58] = 16'd1528;
        rom[ 59] = 16'd1574;
        rom[ 60] = 16'd1622;
        rom[ 61] = 16'd1672;
        rom[ 62] = 16'd1723;
        rom[ 63] = 16'd1776;
        rom[ 64] = 16'd1892;   // exp(2.0)*256 = 1892
        rom[ 65] = 16'd1950;
        rom[ 66] = 16'd2010;
        rom[ 67] = 16'd2072;
        rom[ 68] = 16'd2135;
        rom[ 69] = 16'd2200;
        rom[ 70] = 16'd2268;
        rom[ 71] = 16'd2337;
        rom[ 72] = 16'd2409;
        rom[ 73] = 16'd2483;
        rom[ 74] = 16'd2559;
        rom[ 75] = 16'd2637;
        rom[ 76] = 16'd2718;
        rom[ 77] = 16'd2801;
        rom[ 78] = 16'd2887;
        rom[ 79] = 16'd2975;
        rom[ 80] = 16'd3066;
        rom[ 81] = 16'd3160;
        rom[ 82] = 16'd3257;
        rom[ 83] = 16'd3357;
        rom[ 84] = 16'd3460;
        rom[ 85] = 16'd3566;
        rom[ 86] = 16'd3675;
        rom[ 87] = 16'd3787;
        rom[ 88] = 16'd3903;
        rom[ 89] = 16'd4023;
        rom[ 90] = 16'd4146;
        rom[ 91] = 16'd4274;
        rom[ 92] = 16'd4405;
        rom[ 93] = 16'd4540;
        rom[ 94] = 16'd4679;
        rom[ 95] = 16'd4823;
        rom[ 96] = 16'd5143;   // exp(3.0)*256 = 5143
        rom[ 97] = 16'd5302;
        rom[ 98] = 16'd5465;
        rom[ 99] = 16'd5634;
        rom[100] = 16'd5807;
        rom[101] = 16'd5986;
        rom[102] = 16'd6170;
        rom[103] = 16'd6359;
        rom[104] = 16'd6554;
        rom[105] = 16'd6755;
        rom[106] = 16'd6962;
        rom[107] = 16'd7175;
        rom[108] = 16'd7395;
        rom[109] = 16'd7622;
        rom[110] = 16'd7856;
        rom[111] = 16'd8097;
        rom[112] = 16'd8346;
        rom[113] = 16'd8603;
        rom[114] = 16'd8868;
        rom[115] = 16'd9141;
        rom[116] = 16'd9423;
        rom[117] = 16'd9713;
        rom[118] = 16'd10013;
        rom[119] = 16'd10323;
        rom[120] = 16'd10642;
        rom[121] = 16'd10971;
        rom[122] = 16'd11311;
        rom[123] = 16'd11661;
        rom[124] = 16'd12023;
        rom[125] = 16'd12397;
        rom[126] = 16'd12782;
        rom[127] = 16'd13181;

        // Negative side (signed -128..-1): exp(signed_i/32)*256
        rom[128] = 16'd5;      // exp(-128/32)*256 = exp(-4)*256 = 4.7
        rom[129] = 16'd5;
        rom[130] = 16'd5;
        rom[131] = 16'd5;
        rom[132] = 16'd5;
        rom[133] = 16'd6;
        rom[134] = 16'd6;
        rom[135] = 16'd6;
        rom[136] = 16'd6;
        rom[137] = 16'd6;
        rom[138] = 16'd7;
        rom[139] = 16'd7;
        rom[140] = 16'd7;
        rom[141] = 16'd7;
        rom[142] = 16'd8;
        rom[143] = 16'd8;
        rom[144] = 16'd8;      // exp(-112/32)*256 = exp(-3.5)*256 ~ 7.7
        rom[145] = 16'd8;
        rom[146] = 16'd9;
        rom[147] = 16'd9;
        rom[148] = 16'd9;
        rom[149] = 16'd10;
        rom[150] = 16'd10;
        rom[151] = 16'd10;
        rom[152] = 16'd11;
        rom[153] = 16'd11;
        rom[154] = 16'd12;
        rom[155] = 16'd12;
        rom[156] = 16'd12;
        rom[157] = 16'd13;
        rom[158] = 16'd13;
        rom[159] = 16'd14;
        rom[160] = 16'd14;     // exp(-96/32)*256 = exp(-3)*256 ~ 12.7
        rom[161] = 16'd15;
        rom[162] = 16'd15;
        rom[163] = 16'd16;
        rom[164] = 16'd16;
        rom[165] = 16'd17;
        rom[166] = 16'd17;
        rom[167] = 16'd18;
        rom[168] = 16'd18;
        rom[169] = 16'd19;
        rom[170] = 16'd20;
        rom[171] = 16'd20;
        rom[172] = 16'd21;
        rom[173] = 16'd22;
        rom[174] = 16'd22;
        rom[175] = 16'd23;
        rom[176] = 16'd24;
        rom[177] = 16'd24;
        rom[178] = 16'd25;
        rom[179] = 16'd26;
        rom[180] = 16'd27;
        rom[181] = 16'd28;
        rom[182] = 16'd28;
        rom[183] = 16'd29;
        rom[184] = 16'd30;
        rom[185] = 16'd31;
        rom[186] = 16'd32;
        rom[187] = 16'd33;
        rom[188] = 16'd34;
        rom[189] = 16'd35;
        rom[190] = 16'd36;
        rom[191] = 16'd37;
        rom[192] = 16'd35;     // exp(-64/32)*256 = exp(-2)*256 ~ 34.6
        rom[193] = 16'd36;
        rom[194] = 16'd37;
        rom[195] = 16'd38;
        rom[196] = 16'd40;
        rom[197] = 16'd41;
        rom[198] = 16'd42;
        rom[199] = 16'd43;
        rom[200] = 16'd45;
        rom[201] = 16'd46;
        rom[202] = 16'd48;
        rom[203] = 16'd49;
        rom[204] = 16'd51;
        rom[205] = 16'd52;
        rom[206] = 16'd54;
        rom[207] = 16'd56;
        rom[208] = 16'd57;
        rom[209] = 16'd59;
        rom[210] = 16'd61;
        rom[211] = 16'd63;
        rom[212] = 16'd65;
        rom[213] = 16'd67;
        rom[214] = 16'd69;
        rom[215] = 16'd71;
        rom[216] = 16'd73;
        rom[217] = 16'd75;
        rom[218] = 16'd78;
        rom[219] = 16'd80;
        rom[220] = 16'd82;
        rom[221] = 16'd85;
        rom[222] = 16'd88;
        rom[223] = 16'd90;
        rom[224] = 16'd94;     // exp(-32/32)*256 = exp(-1)*256 ~ 94
        rom[225] = 16'd97;
        rom[226] = 16'd100;
        rom[227] = 16'd103;
        rom[228] = 16'd106;
        rom[229] = 16'd110;
        rom[230] = 16'd113;
        rom[231] = 16'd116;
        rom[232] = 16'd120;
        rom[233] = 16'd124;
        rom[234] = 16'd127;
        rom[235] = 16'd131;
        rom[236] = 16'd135;
        rom[237] = 16'd139;
        rom[238] = 16'd144;
        rom[239] = 16'd148;
        rom[240] = 16'd153;    // exp(-16/32)*256 = exp(-0.5)*256 ~ 155
        rom[241] = 16'd158;
        rom[242] = 16'd162;
        rom[243] = 16'd167;
        rom[244] = 16'd172;
        rom[245] = 16'd178;
        rom[246] = 16'd183;
        rom[247] = 16'd189;
        rom[248] = 16'd195;
        rom[249] = 16'd201;
        rom[250] = 16'd207;
        rom[251] = 16'd213;
        rom[252] = 16'd220;
        rom[253] = 16'd227;
        rom[254] = 16'd234;
        rom[255] = 16'd241;    // exp(-1/32)*256 ~ 248
    end

    // ----------------------------------------------------------------
    // Registered read (1-cycle latency)
    // ----------------------------------------------------------------
    always_ff @(posedge clk) begin
        data_out <= rom[addr];
    end

endmodule
